//Data memory module --Rishi
module dataMemory(
input wire CLK,
input wire [31:0] ALUResult,
input wire [31:0] WriteData,
input wire WE,



);
